`define num_of_txns 20
